hello whats good
  
